library verilog;
use verilog.vl_types.all;
entity CLA_adder64bit_tb is
end CLA_adder64bit_tb;
