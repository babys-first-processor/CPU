library verilog;
use verilog.vl_types.all;
entity dff_async_reset_tb is
end dff_async_reset_tb;
