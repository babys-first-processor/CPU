library verilog;
use verilog.vl_types.all;
entity tribuf_tb is
end tribuf_tb;
