module rom_case(out, address);
output reg[31:0] out;
input [11:0] address;


always @*
	begin
			case (address)
				12'h800: out <= 32'b1001000100_000000000000_11111_00000;
				12'h801: out <= 32'b1001000100_000000000001_11111_00001;
				12'h802: out <= 32'b10001011000_00000_000000_00001_00010;
				12'h803: out <= 32'b10001011000_11111_000000_00001_00000;
				12'h804: out <= 32'b10001011000_11111_000000_00010_00001;
				12'h805: out <= 32'b1111000100_111111111111_00000_11111;
				12'h806: out <= 32'b01010100_0000000100000000000_0_1100;
				12'h807: out <= 32'b000101_00000000000000100000000010;
				//...
				12'h8FD: out <= 32'b00000000111111110000000011111111;
				12'h8FE: out <= 32'b11111111000000001111111100000000;
				12'h8FF: out <= 32'b11111111111111111111111111111111;
				default: out <= 32'b00000000000000000000000000000000;
				//this should be updated eventually to use .mem files from assembler?
			endcase
	end
endmodule

			