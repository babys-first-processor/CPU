library verilog;
use verilog.vl_types.all;
entity regfile32x64_tb is
end regfile32x64_tb;
